`define ADDRESS_SIZE                64
`define BLOCK_SIZE                  64
`define BUS_DATA_WIDTH              64
`define BUS_TAG_WIDTH               13
`define DATA_SIZE                   64
`define DIRTY                       1
`define IMMEDIATE_SIZE              64
`define INDEX_SIZE                  32 
`define INDEX_SIZE_B                $clog2(`INDEX_SIZE - 1)
`define INDEXES_PER_WAY             32
`define INSTRUCTION_SIZE            32
`define LSQ_SIZE                    1
`define MEM_READ                    0'h1100
`define NUMBER_OF_REGISTERS         32
`define NUMBER_OF_REGISTERS_B       $clog2(`NUMBER_OF_REGISTERS - 1)
`define OFFSET_SIZE                 64 
`define OFFSET_SIZE_B               $clog2(`OFFSET_SIZE - 1)
`define CELLS_NEEDED                8
`define CELLS_NEEDED_B              $clog2(`CELLS_NEEDED - 1)
`define ROB_SIZE                    `LSQ_SIZE
`define RS_SIZE                     `ROB_SIZE
`define TAG_SIZE_B                  64 - (`OFFSET_SIZE_B + `INDEX_SIZE_B)
`define VALID                       1
`define WAYS                        4
`define WAYS_B                      $clog2(`WAYS - 1)


// Data Structure Lengths
`define CONTROL_BITS_SIZE           $bits(control_bits)



// OFFSET bits will alawys be a multiple of 4
// TAG SIZE + INDEX + OFFSET
//   53         5       6

typedef logic [`TAG_SIZE_B - 1 : 0] cache_tag; 
typedef logic [`INDEX_SIZE_B - 1 : 0] cache_index;
typedef logic [`OFFSET_SIZE_B - 1 : 0] cache_offset;
// CACHE CONSTANTS
typedef struct packed {
  cache_tag tag;
  cache_index index;
  cache_offset offset;
} cache_address;

// Cache Block
// Block size = 32 * (1 + 1 + 53 + 3 * 64) = 18176 bits
typedef logic [`DATA_SIZE - 1 : 0] cache_cell; // One Cell of Size 64
typedef struct packed {
  logic valid;
  logic dirty;
  logic [`TAG_SIZE_B - 1 : 0] tag;
  cache_cell [`CELLS_NEEDED - 1 : 0] cache_cells; // 64 byte offset (8 cells)
} cache_line;
typedef cache_line[`INDEXES_PER_WAY - 1 : 0] cache_block;
typedef cache_block [`WAYS - 1 : 0] full_cache;








// Memory Instruction Type
typedef enum logic[3:0] { 
        LB, LBU, LH, LHU, LW, LWU, LD,
        SB, SH, SW, SD 
      } memory_instruction_type;

// ALU operation
typedef enum logic [5:0] {
  // Normal ALU
  ADD, SUB, AND, OR, XOR,
  SLT, SRL, SRA, SLL,
  ADDW, SUBW, SLTW, SRAW, SRLW, SLLW,
  BEQ, BNE, BGE, BLT, BGEU, BLTU,
  //M extention
  MUL, MULH, MULSU, MULHU, MULHSU,
  MULW, DIV, DIVU, REM,
  REMU, DIVW, DIVUW,
  REMW, REMUW
} alu_operation;

typedef struct packed {
  logic alusrc;                       // ALU source (rs2 or imm)
  logic apc;                          // Adding PC
  logic cjump;                        // Conditional Jump
  logic ecall;                        // e-call
  logic memtoreg;                     // Memory To Register
  logic memwr;                        // Memory Write
  logic regwr;                        // Register Write
  logic ucjump;                       // Unconditional Jump
  logic unsupported;                  // *Unsuppored Instruction
  logic usign;                        // Unsigned
  alu_operation aluop;                // ALU Operation
  memory_instruction_type memorytype; // Memory Instruction Type
} control_bits;









/////////////////////////////////////////////////////////////////////////////////
/********************************** REGISTERS **********************************/
/////////////////////////////////////////////////////////////////////////////////
// Register between fetch and decode
typedef struct packed {
  logic [`INSTRUCTION_SIZE - 1 : 0] instruction;
} fetch_decode_register;

// Register between decode and register fetch
typedef struct packed {
  logic [`INSTRUCTION_SIZE - 1 : 0] instruction;
	logic [`NUMBER_OF_REGISTERS_B - 1 : 0] rs1;
  logic [`NUMBER_OF_REGISTERS_B - 1 : 0] rs2;
  logic [`NUMBER_OF_REGISTERS_B - 1 : 0] rd;
	logic [`IMMEDIATE_SIZE - 1 : 0] imm;
	logic [`CONTROL_BITS_SIZE - 1 : 0] ctrl_bits;
} decode_registers_register;

// Register between register fetch and dipatch
typedef struct packed {
  logic [`INSTRUCTION_SIZE - 1 : 0] instruction;
	logic [`NUMBER_OF_REGISTERS_B - 1 : 0] rs1;
  logic [`NUMBER_OF_REGISTERS_B - 1 : 0] rs2;
  logic [`NUMBER_OF_REGISTERS_B - 1 : 0] rd;
  logic [`DATA_SIZE - 1 : 0] rs1_value;
  logic [`DATA_SIZE - 1 : 0] rs2_value;
	logic [`IMMEDIATE_SIZE - 1 : 0] imm;
	logic [`CONTROL_BITS_SIZE - 1 : 0] ctrl_bits;
} registers_dispatch_register;



/////////////////////////////////////////////////////////////////////////////////
/********************************** HARDWARE ***********************************/
/////////////////////////////////////////////////////////////////////////////////
typedef struct packed {
  logic in_rob;
  int tag;
} map_table_entry;

typedef struct packed {
  logic ready
  int tag;
  logic [`NUMBER_OF_REGISTERS_B - 1 : 0] register_destination;
  logic [`DATA_SIZE - 1 : 0] value;
  control_bits ctrl_bits;
} rob_entry;

typedef struct packed {
  logic busy;
  int id;
  int tag;
  int tag_1;
  int tag_2;
  logic [`DATA_SIZE - 1 : 0] value_1;
  logic [`DATA_SIZE - 1 : 0] value_2;
  control_bits ctrl_bits;
} rs_entry;

typedef struct packed {
  memory_instruction_category category;
  memory_instruction_type memory_type;
  int tag;
  logic [`ADDRESS_SIZE - 1 : 0] address;
  logic [`DATA_SIZE - 1 : 0] value;
} lsq_entry;


