`include "Sysbus.defs"
`include "src/consts.sv"
`include "src/cache.sv"

module top
#(
  BUS_DATA_WIDTH = 64,
  BUS_TAG_WIDTH = 13
)
(
  input  clk,
         reset,

  // 64-bit addresses of the program entry point and initial stack pointer
  input  [63:0] entry,
  input  [63:0] stackptr,
  input  [63:0] satp,
  
  // interface to connect to the bus
  output bus_reqcyc,
  output bus_respack,
  output [BUS_DATA_WIDTH-1:0] bus_req,
  output [BUS_TAG_WIDTH-1:0] bus_reqtag,
  input  bus_respcyc,
  input  bus_reqack,
  input  [BUS_DATA_WIDTH-1:0] bus_resp,
  input  [BUS_TAG_WIDTH-1:0] bus_resptag
);

  logic [63:0] pc;

  always @ (posedge clk)
    if (reset) begin
      pc <= entry;
    end else begin
      $display("Hello World!  @ %x", pc);
      $finish;
    end

  initial begin
    $display("Initializing top, entry point = 0x%x", entry);
  end
endmodule
